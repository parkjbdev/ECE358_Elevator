`timescale 100ms / 100ms

module controller(
  input clk,
  input set_clk,
  input [2:0] src_input,
  input [2:0] dest_input,
  input direction_input, // up = 1, down = 0
  output [2:0] ev_floor
);
  reg [2:0] target_floor_input;
  wire ev_door;

  mover u_mover(
    // inputs
    .dest_input(target_floor_input),
    // outputs
    .ev_floor_output(ev_floor),
    .ev_door_output(ev_door)
  );

  // Input Saving Registers
  reg [2:0] src1_input, src2_input;
  reg [2:0] dest1_input, dest2_input;
  reg direction1_input, direction2_input;

  // Variables
  reg [1:0] done, on_board;

  initial begin
    done = 2'b11;
    on_board = 2'b00;
  end

  // Assigning Inputs
  always @(posedge set_clk) begin
    // Assertion
    if (src_input == dest_input)
      $display("Input Assertion Failed");
    else if (src_input > dest_input & direction_input == 1)
      $display("Input Assertion Failed");
    else if (src_input < dest_input & direction_input == 0)
      $display("Input Assertion Failed");
    else begin
      casex (done)
        2'b00: $display("Elevator busy");
        2'bx1: begin
          $display("1 is assigned");
          done = done & 2'b10; // #1 is not done
          src1_input = src_input;
          dest1_input = dest_input;
          direction1_input = direction_input;
        end
        2'b1x: begin
          $display("2 is assigned");
          done = done & 2'b01; // #2 is not done
          src2_input = src_input;
          dest2_input = dest_input;
          direction2_input = direction_input;
        end
      endcase
    end
  end

  // Only when elevator door opens
  always @(posedge ev_door) begin
    // On Destination Arrival
    // 1st person
    // done: 2'bx0, on_board: 2'bx0
    if ((done == 2'b10 | done == 2'b00) & (on_board == 2'b10 | on_board == 2'b00) & ev_floor == src1_input) // If 1st rides
    begin
      target_floor_input = src1_input; // open and close door
      on_board = on_board + 2'b01; // on_board = 2'bx1;
    end
    // done: 2'bx0, on_board: 2'bx1
    else if ((done == 2'b10 | done == 2'b00) & (on_board == 2'b11 | on_board == 2'b01) & ev_floor == dest1_input) // If 1st person arrived dest.
    begin
      target_floor_input = dest1_input; // open and close door
      done = done + 2'b01; // done = 2'bx1
      on_board = on_board & 2'b10; // on_board = 2'bx0;
    end

    // 2nd person
    // done: 2'b0x, on_board: 2'b0x
    if ((done == 2'b01 | done == 2'b00) & (on_board == 2'b01 | on_board == 2'b00) & ev_floor == src2_input) // If 2nd rides
    begin
      target_floor_input = src2_input; // open and close door
      on_board = on_board + 2'b10; // on_board = 2'b1x;
    end
    // done: 2'b0x, on_board: 2'b1x
    else if ((done == 2'b01 | done == 2'b00) & (on_board == 2'b10 | on_board == 2'b11) & ev_floor == dest2_input) // If 2nd person arrived dest.
    begin
      target_floor_input = dest2_input; // open and close door
      done = done + 2'b10; // done = 2'b1x
      on_board = on_board & 2'b01; // on_board = 2'b0x;
    end
  end

  always @(clk) begin
    if (done == 2'b00)
    begin
      if (direction1_input == 1 & direction2_input == 1)
      begin
        if (on_board == 2'b01) // only 1 is on ride
        begin
          if (src2_input > ev_floor)
          begin
            if (src2_input < dest1_input) target_floor_input = src2_input;
            else target_floor_input = dest1_input;
          end
        end

        else if (on_board == 2'b10) // only 2 is on ride
        begin
          if (src1_input > ev_floor)
          begin
            if (src1_input < dest2_input) target_floor_input = src1_input;
            else target_floor_input = dest2_input;
          end
        end

        else if (on_board == 2'b00) // 1 and 2 both is not on ride yet
        begin
          if (src1_input < src2_input) target_floor_input = src1_input;
          else target_floor_input = src2_input;
        end
  
        else if (on_board == 2'b11) // 1 and 2 is both on ride
        begin
          if (dest1_input < dest2_input) target_floor_input = dest1_input;
          else target_floor_input = dest2_input;
        end
      end

      else if (direction1_input == 0 & direction2_input == 0)
      begin
        if (on_board == 2'b01) // only 1 is on ride
        begin
          if (src2_input < ev_floor)
          begin
            if (src2_input > dest1_input) target_floor_input = src2_input;
            else target_floor_input = dest1_input;
          end
        end

        else if (on_board == 2'b10) // only 2 is on ride
        begin
          if (src1_input < ev_floor)
          begin
            if (src1_input > dest2_input) target_floor_input = src1_input;
            else target_floor_input = dest2_input;
          end
        end

        else if (on_board == 2'b00) // 1 and 2 both is not on ride yet
        begin
          if (src1_input > src2_input) target_floor_input = src1_input;
          else target_floor_input = src2_input;
        end
  
        else if (on_board == 2'b11) // 1 and 2 is both on ride
        begin
          if (dest1_input > dest2_input) target_floor_input = dest1_input;
          else target_floor_input = dest2_input;
        end
      end
      else
      begin
        if (on_board == 2'b00) target_floor_input = src1_input;
        else if (on_board == 2'b01) target_floor_input = dest1_input;
      end
    end
    else if (done == 2'b10) // 1 is not done
    begin
      if (on_board == 2'b00 | on_board == 2'b10) target_floor_input = src1_input;
      else if (on_board == 2'b01 | on_board == 2'b11) target_floor_input = dest1_input;
    end
    else if (done == 2'b01) // 2 is not done
    begin
      if (on_board == 2'b00 | on_board == 2'b01) target_floor_input = src2_input;
      else if (on_board == 2'b10 | on_board == 2'b11) target_floor_input = dest2_input;
    end
  end


  // Output
  // assign current_floor_output = ev_floor;
endmodule

module mover(
  input[2:0] dest_input,
  output[2:0] ev_floor_output,
  output ev_door_output
);

reg clk;
initial clk = 0;
always #1 clk = ~clk;

// States
parameter IDLE_OPENED = 2'b11;
parameter IDLE_CLOSED = 2'b00;
parameter MOVING_UP = 2'b01;
parameter MOVING_DOWN = 2'b10;

// State
reg[1:0] state;
initial state = IDLE_CLOSED;

// Arrival Flag
reg arrived;
initial arrived = 1;

always @(ev_floor or dest_input or ev_door)
  case (state)
    IDLE_CLOSED:
    begin
      if (dest_input > ev_floor_output) state = MOVING_UP;
      else if (dest_input < ev_floor_output) state = MOVING_DOWN;
      else if (arrived == 0) state = IDLE_OPENED;
      else state = IDLE_CLOSED;
    end

    IDLE_OPENED:
    begin
      if (arrived == 1) state = IDLE_CLOSED;
      arrived = 1;
    end

    MOVING_DOWN:
    begin
      arrived = 0;
      if (dest_input < ev_floor_output) state = MOVING_DOWN;
      else state = IDLE_CLOSED;
    end

    MOVING_UP:
    begin
      arrived = 0;
      if (dest_input > ev_floor_output) state = MOVING_UP;
      else state = IDLE_CLOSED;
    end
 
    default: state = IDLE_CLOSED;
  endcase

// Elevator Module
reg ev_door_open;
reg [1:0] ev_updown;
wire ev_door;
wire [2:0] ev_floor;


elevator u_elevator(
  .clk(clk),
  // inputs
  .door_open(ev_door_open),
  .updown(ev_updown),
  // outputs
  .door(ev_door),
  .floor(ev_floor)
);

always @(state) begin
  case (state)
    IDLE_CLOSED:
    begin
      ev_door_open = 0;
      ev_updown = 2'b00;
    end

    IDLE_OPENED:
    begin
      // arrived = 1;
      ev_door_open = 1;
      ev_updown = 2'b00;
    end

    MOVING_DOWN:
    begin
      // arrived = 0;
      ev_door_open = 0;
      ev_updown = 2'b10;
    end

    MOVING_UP:
    begin
      // arrived = 0;
      ev_door_open = 0;
      ev_updown = 2'b01;
    end

    default:
    begin
      // arrived = 1;
      ev_door_open = 0;
      ev_updown = 2'b00;
    end
  endcase
end

assign ev_floor_output = ev_floor;
assign ev_door_output = ev_door;

endmodule
